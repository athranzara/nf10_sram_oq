`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   19:10:55 02/16/2015
// Design Name:   Axi2Fifo_asyn
// Module Name:   /local/scratch/jz377/git_repo/nf10_sram_oq/pcores/nf10_sram_output_queue_v1_00_a/hdl/verilog/axi2fifo_asyn_tb.v
// Project Name:  nf10_sram_output_queue
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: Axi2Fifo_asyn
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module axi2fifo_asyn_tb;

	// Inputs
	reg clk;
	reg reset;
	reg memclk;
	reg memreset;
	reg tvalid;
	reg [255:0] tdata;
	reg [31:0] tstrb;
	reg [127:0] tuser;
	reg tlast;
	reg output_enable;

	// Outputs
	wire tready;
	wire [201:0] dout;
	wire dout_valid;
	wire [4:0] oq;

	// Instantiate the Unit Under Test (UUT)
	Axi2Fifo_asyn uut (
		.clk(clk), 
		.reset(reset), 
		.memclk(memclk), 
		.memreset(memreset), 
		.tvalid(tvalid), 
		.tready(tready), 
		.tdata(tdata), 
		.tstrb(tstrb), 
		.tuser(tuser), 
		.tlast(tlast), 
		.dout(dout), 
		.dout_valid(dout_valid), 
		.output_enable(output_enable), 
		.oq(oq)
	);
	
	
localparam [95:0]   tuser_para1 = 96'b0;
localparam [7:0]    tuser_para2 = 8'b10101111;
localparam [23:0]   tuser_para3 = 24'b1;
localparam [7:0]    tuser_para2_2 = 8'b11101010;

reg [7:0]   i;
reg [255:0] tdata1;
reg [255:0] tdata2;
reg         packet_num;
reg [1:0]   axis_state,next_axis_state;

localparam PACKET_LEN = 20;
localparam GETREADY = 0;
localparam TRANSMISSION = 1;

reg [255:0] next_tdata;
reg [127:0] next_tuser;
reg [31:0]  next_tstrb;
reg         next_tvalid;

/* axis simulator*/
//always @ (posedge clk) begin
//    if (reset) begin
//        axis_state <= 0;
//        tdata <= {256{1'b0}};
//        tuser <= {128{1'b0}};
//        tstrb <= {32{1'b0}};
//        tvalid<= 1'b0;
//    end
//    else begin
//        axis_state <= next_axis_state;
//        tdata <= next_tdata;
//        tuser <= next_tuser;
//        tstrb <= next_tstrb;
//        tvalid<= next_tvalid;
//    end
//end

//always @ * begin
//next_axis_state = axis_state;
//next_tdata = tdata;
//next_tuser = tuser;
//next_tstrb = tstrb;
//next_tvalid = tvalid;

//end

always @ * begin
    if (reset) begin
        axis_state = 0;
        next_axis_state = 0;
    end
    else begin
        axis_state = next_axis_state;
    end

end

    always @ * begin
        tlast = 1'b0;
        tstrb = tstrb;
        if (i == PACKET_LEN) begin
            tlast = 1'b1;
            tstrb = 32'h000fffff;
        end

    end

//always @ * begin
//    next_axis_state = 
//end

always @ (posedge clk) begin
    case (axis_state)
    GETREADY:       begin
                        if (~reset) begin
                            if (packet_num == 0) begin
                                tdata <= tdata1;
                                tuser <= {tuser_para1,tuser_para2,tuser_para3};
                                tvalid <= 1'b1;
                                tstrb <= 32'hffffffff;
                                packet_num <= 1;
                                i = 0;
                            end
                            else if (packet_num == 1) begin
                                tstrb <= 32'hffffffff;
                                tdata <= tdata2;
                                tuser <= {tuser_para1,tuser_para2_2,tuser_para3};
                                tvalid <= 1'b1;
                                packet_num <=0;
                                i = 0;
                            end
                            next_axis_state <= TRANSMISSION;
                        end
                        

                    end
    
    TRANSMISSION:   begin
                        if (tlast) begin
                            next_axis_state <= GETREADY;
                        end
                        else if (tready) begin
                        tdata <= tdata + 256'd1;
                        i = i + 1;
                        end
                    end
                    
    default:        begin
                    tvalid <= 0;
                    tdata <= 256'bz;
                    tuser <= 128'bz;
                    tstrb <= 32'bz;
                    /*pause*/
                    end
    endcase
    
    

end

/* end of axis simulator*/

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		memclk = 0;
		memreset = 1;
		tvalid = 0;
		tdata = 0;
		tdata1 = 50;
		tdata2 = 200;
		tstrb = 0;
		tuser = 0;
		output_enable = 0;
		i = 0;
		packet_num = 0;

		// Wait 100 ns for global reset to finish
		#20;
        reset = 1'b0;
        memreset = 1'b0;
		// Add stimulus here
		output_enable = 1'b1;


	end
	
    always #3.125   begin
        clk = ~clk;         // 160MHz
    end
    

    always #2 begin
        memclk = ~memclk;   // 250MHz
    end
    
// simulatre arbitor behavior

always @ (posedge memclk) begin
    
end
    
    
      
endmodule

